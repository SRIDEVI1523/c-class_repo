// Copyright (c) 2020 IIT Madras. see LICENSE.iitm for more details on licensing terms
/*
Author: Neel Gala, neelgala@incoresemi.com
Created on: Monday 21 June 2021 09:07:59 PM

*/
/*doc:overview:
This is the write-back stage of the pipeline where all instructions retire. By the time an
instructino reaches this stage it has been narrowed down via some of the previous stages into one of
the following categories of operations that can be performed in this stage:

  - SYSTEM: either xRET operations or CSR access operations.
  - TRAP: The instruction has encountered a trap during its operation in one of the previous stages.
  - BASEOUT: The instruction retirement includes a simple update to the registerfile
  - MEMOP: The instruction is either a cached store/atomic operation or an non-cached/IO memory op.

Each of the above have a unique ISB feeding in respective instructions to this module. This module
uses the fuid from the previous stage,  which maintains the order of instructions to find out which
ISB must be polled for the retiring/committing the next instruction.

Operations which can take multiple cycles in this stage are : CSR operations if daisy-chain is more
than 1 level deep; IO/non-cached Memory Operations may also take significantly longer in this stage
to complete.

All other ops will take a single cycle to complete.

When in simulation mode, this module will offload the commit-log packet to the test-bench via a
single Default-Reg (DReg) interface.

This module also instantiates the csrbox module, which hosts all the csrs and also the routines to
perform a trap or an xRet operation. Certain csr interfaces are simply bypassed along this module so
that they are exposed at the next hiegher level to rest of the pipeline and design.

*/
package stage5 ;

import FIFOF        :: * ;
import Vector       :: * ;
import SpecialFIFOs :: * ;
import FIFOF        :: * ;
import TxRx         :: * ;
import DefaultValue :: * ;
import Assert       :: * ;
import Connectable  :: * ;

`include "Logger.bsv"
`include "trap.defines"

import pipe_ifcs    :: * ;
import dcache_types :: * ;
import csrbox       :: * ;
import csr_types    :: * ;
import ccore_types  :: * ;
import DReg         :: * ;


interface Ifc_stage5;
`ifdef debug
  interface Ifc_s5_debug debug;
`endif
`ifdef perfmonitors
  interface Ifc_s5_perfmonitors perf;
`endif
  interface Ifc_s5_rx rx;
  interface Ifc_s5_interrupts interrupts;
  interface Ifc_s5_common common;
  interface Ifc_s5_cache cache;
  interface Ifc_s5_csrs csrs;
endinterface:Ifc_stage5

`ifdef stage5_noinline
/*doc:module: */
(*synthesize*)
`endif
`ifdef simulate
(*preempts = "rl_writeback_memop, rl_no_op"*)
(*preempts = "rl_writeback_trap, rl_no_op"*)
(*preempts = "rl_writeback_system, rl_no_op"*)
(*preempts = "rl_writeback_baseout, rl_no_op"*)
`endif
module mkstage5#(parameter Bit#(`xlen) hartid) (Ifc_stage5);

  /*doc:submodules: The following instantiates all the RX virtual fifos*/
  RX#(SystemOut) rx_systemout <- mkRX;
  RX#(TrapOut)   rx_trapout <- mkRX;
  RX#(BaseOut)   rx_baseout <- mkRX;
  RX#(WBMemop)   rx_memio <- mkRX;
  RX#(CUid)      rx_fuid <- mkRX;
`ifdef rtldump
  RX#(CommitLogPacket) rx_commitlog <- mkRX;
`endif
 
  /*doc:submodules: The following instantiates the csr module generated by csrbox*/
  Ifc_csrbox csr <- mk_csrbox();

  /*doc:reg: This register holds the local epoch value of this stage*/
  Reg#(Bit#(1)) rg_epoch <- mkReg(0);

  /*doc:reg: This register when set is used to indicate that we need wait for the csrbox to respond*/
  Reg#(Bool) rg_csr_wait <- mkReg(False);

  /*doc:wire wire that carries the commit data that needs to be written to the integer register
   * file. IN cases of traps and instructions that need to be dropped, writing to this wire can be
   * used to release the lock on a register in the score-board*/
  Wire#(CommitData) wr_commit <- mkWire();

  /*doc:wire: This wire is used to indicate the rest of the pipeline that this stage has generated a
  * flush. In case of post-fenceI/sfence this signal also holds fields which are used to indicate
  * the I$ about a possible fenceI or sfence on the ITLB*/
  Wire#(WBFlush) wr_flush <- mkDWire(defaultValue);

  /*doc:wire: When set to True causes an increment in the minstret counter. Note in case of a csr
  * operation that writes a value to minstret. The new value of minstret at the end of the cycle
  * would be write-value + 1.*/
  Wire#(Bool) wr_increment_minstret <- mkDWire(False);

  /*doc:reg: This register when set indicates that an IO memory operation is in progress*/
  Reg#(Bool) rg_ioop_init <- mkReg(False);

  /*doc:wire: This wire holds the response of an IO memory operation */
  Wire#(Maybe#(DMem_core_response#(TMul#(`dwords,8),`desize))) wr_ioop_response <- mkDWire(tagged Invalid);

  /*doc:wire: this wire holds the epoch value of the IO memory store/atomic operation that is
   * waiting to be committed/dropped. Writing a value to this wire triggers an IO operation*/
  Wire#(Bit#(1)) wr_commit_ioop <- mkWire();

`ifdef dcache
  /*doc:wire: this wire holds the epoch value of the cached memory store/atomic operation that is
   * waiting to be committed/dropped*/
  Wire#(Tuple2#(Bit#(1), Bit#(TLog#(`dsbsize)))) wr_commit_cacheop <- mkWire();
`endif    
`ifdef debug
  /*doc:submodules: connection back to the csrs to stop counters*/
  mkConnection(csr.ma_stop_count, csr.mv_stop_count);
`endif
`ifdef rtldump
  /*doc:reg: When an instruction commits, this register holds the commit log packet in the next
   * cycle which can be consumed by the test-bench to write into a file*/
  Reg#(Maybe#(CommitLogPacket)) rg_commitlog <- mkDReg(tagged Invalid);
`endif
`ifdef perfmonitors
  /*doc:wire: wire to increment when exceptions detected*/
  Wire#(Bit#(1)) wr_count_exceptions <- mkDWire(0);
  /*doc:wire: wire to increment when interrupts detected*/
  Wire#(Bit#(1)) wr_count_interrupts <- mkDWire(0);
  /*doc:wire: wire to increment when csr-ops detected*/
  Wire#(Bit#(1)) wr_count_csrops <- mkDWire(0);
  /*doc:wire: wire to increment when micro-traps are detected*/
  Wire#(Bit#(1)) wr_count_microtrap <- mkDWire(0);
`endif

  let csr_response = csr.mv_core_resp;
  let epochs_match = rg_epoch == rx_fuid.u.first.epochs;

`ifdef simulate
  rule rl_no_op;
    `logLevel( stage5, 0, $format("[%2d]STAGE5: No Instr to commit", hartid))
  endrule: rl_no_op
`endif

  /*doc:rule: This rule handles all traps there were detected/raised in any of the previous stages
  * for any given instruction. The rule also checks if the micro-trap is generated and acts
  * accordingly. For a regular trap like load-access/load-page-fault, the load instruction would
  * have locked a register in the score-board and would thus require to be released inspite of
  * taking of the fault. To ensure this release, we update the wr_commit signal to make this release
  * on the destination register*/
  rule rl_writeback_trap(rx_fuid.u.first.insttype == TRAP );
    let trapout = rx_trapout.u.first;
    let fuid = rx_fuid.u.first;
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : PC:%h",hartid,fuid.pc))
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : Trap: ",hartid, fshow(trapout)))
    wr_commit <= CommitData{addr: fuid.rd, data: ?, unlock_only:True
                          `ifdef no_wawstalls , id: fuid.id `endif
                           `ifdef spfpu rdtype: fuid.rdtype `endif };

    if (epochs_match) begin
    `ifdef microtrap_support
      if (trapout.is_microtrap) begin
        if (trapout.cause == `Sfence_rerun || trapout.cause == `FenceI_rerun || 
            trapout.cause == `CSR_rerun 
					`ifdef hypervisor || trapout.cause == `Hfence_rerun `endif ) begin
          let _fencei = (trapout.cause == `FenceI_rerun);
          let _sfence = (trapout.cause == `Sfence_rerun);
  			  let _hfence = (trapout.cause == `Hfence_rerun);
          wr_flush <= WBFlush{flush: True, newpc : fuid.pc , fencei: _fencei 
              `ifdef supervisor , sfence: _sfence `endif 
              `ifdef hypervisor , hfence: _hfence `endif };
          `logLevel( stage5, 0, $format("[%2d]STAGE5 : Redirect PC:%h",hartid, fuid.pc))
        `ifdef perfmonitors
          wr_count_microtrap <= 1;
        `endif
        end
        else begin
          dynamicAssert(False, "Received unexpected Micro-Trap cause");
        end
      end
      else `endif begin
        let tvec <- csr.mav_upd_on_trap(trapout.cause, fuid.pc, trapout.mtval, trapout.mtval2);
        wr_flush <= WBFlush{flush: True, newpc : tvec, fencei: False 
            `ifdef supervisor , sfence: False `endif 
            `ifdef hypervisor , hfence: False `endif };
      `ifdef perfmonitors
        Bit#(1) cause_type = truncateLSB(trapout.cause);
        if (cause_type == 1)
          wr_count_interrupts <= 1;
        else
          wr_count_exceptions <= 1;
      `endif
        `logLevel( stage5, 0, $format("[%2d]STAGE5 : Going to *TVEC:%h",hartid, tvec))
      end
        rx_trapout.u.deq;
        rx_fuid.u.deq;
        rg_epoch <= ~rg_epoch;
      `ifdef rtldump
        rx_commitlog.u.deq;
      `endif
    end
    else begin
      `logLevel( stage5, 0, $format("[%2d]STAGE5 : Dropping instruction",hartid))
      rx_trapout.u.deq;
      rx_fuid.u.deq;
    `ifdef rtldump
      rx_commitlog.u.deq;
    `endif
    end
  endrule:rl_writeback_trap

  /*doc:rule: This rule is used to commit system operations which could be xRET ops or CSR ops.
  * Committing a xRET ops causes a flush to be raised with a new pc coming from the csrbox. In case
  * of CSR ops, one might have to wait for multiple cycles for the execution to complete and then
  * commit the value.*/
  rule rl_writeback_system(rx_fuid.u.first.insttype == SYSTEM ) ;
    let systemout = rx_systemout.u.first;
    let fuid = rx_fuid.u.first;
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : PC:%h",hartid,fuid.pc))
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : ",hartid, fshow(systemout)))
    Bool exit = False;
    if (epochs_match) begin
      if (systemout.funct3 == 0 ) begin // URET, SRET, MRET
        let epc <- csr.mav_upd_on_ret(truncateLSB(systemout.csr_address));
        exit = True;
        wr_flush <= WBFlush{flush: True, newpc : epc, fencei: False
          `ifdef supervisor , sfence: False `endif 
          `ifdef hypervisor , hfence: False `endif };
        rg_epoch <= ~rg_epoch;
          `logLevel( stage5, 0, $format("[%2d]STAGE5 : Redirect PC:%h",hartid,epc))
      end
      else if (!rg_csr_wait) begin
        csr.ma_core_req(CSRReq{csr_address: systemout.csr_address, writedata: systemout.rs1_imm,
            funct3: truncate(systemout.funct3) `ifdef compressed , pc_1: fuid.pc[1] `endif });
      end
  
      if ((systemout.funct3 !=0 && csr_response.hit) || (systemout.funct3==0)) begin
        rg_csr_wait <= False;
        exit = True;
      end
      else begin
        rg_csr_wait <= True;
        `logLevel( stage5, 0, $format("[%2d]STAGE5 : Waiting for CSR-response",hartid))
      end
  
      if (exit) begin
        wr_increment_minstret <= True;
        wr_commit <= CommitData{addr: fuid.rd, data: zeroExtend(csr_response.data), unlock_only:False
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu rdtype: fuid.rdtype `endif };
        rx_systemout.u.deq;
        rx_fuid.u.deq;
      `ifdef perfmonitors
        if (systemout.funct3 != 0)
          wr_count_csrops <= 1;
      `endif
      `ifdef rtldump
        let clogpkt = rx_commitlog.u.first;
        CommitLogCSR _pkt = ?;
        if (clogpkt.inst_type matches tagged CSR .pcsr)
          _pkt = pcsr;
        if (systemout.funct3 == 0) begin
          _pkt.csr_address = 'h300;
          _pkt.wdata = csr.sbread.mv_csr_mstatus;
        end
        _pkt.rdata = csr_response.data;
        clogpkt.inst_type = tagged CSR _pkt;
        clogpkt.mode = csr.mv_prv;
			`ifdef hypervisor
				clogpkt.v = csr.mv_virtual;
			`endif
        rg_commitlog <= tagged Valid clogpkt;
        rx_commitlog.u.deq;
      `endif
      end
    end
    else begin
      `logLevel( stage5, 0, $format("[%2d]STAGE5 : Dropping instruction",hartid))
      wr_commit <= CommitData{addr: fuid.rd, data: ?, unlock_only:True
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu rdtype: fuid.rdtype `endif };
      rx_systemout.u.deq;
      rx_fuid.u.deq;
    `ifdef rtldump
      rx_commitlog.u.deq;
    `endif
    end
  endrule:rl_writeback_system

  /*doc:rule: This rule basically commits regular ops which update the register file. Note that even
  * Loads will land up here. So the commit log packet is not touched since it would be tagged
  * CommitLogMem for Loads which has to be passed on as is to the test-bench*/
  rule rl_writeback_baseout(rx_fuid.u.first.insttype == BASE);
    let fuid = rx_fuid.u.first;
    let baseout = rx_baseout.u.first;
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : PC:%h",hartid,rx_fuid.u.first.pc))
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : Base Op ",hartid, fshow(baseout)))
    if (epochs_match) begin
      wr_increment_minstret <= True;
      `ifdef spfpu csr.ma_set_fflags(baseout.fflags); `endif
      wr_commit <= CommitData{addr: fuid.rd, data: zeroExtend(baseout.rdvalue), unlock_only:False
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu rdtype: fuid.rdtype `endif };
      rx_fuid.u.deq;
      rx_baseout.u.deq;
    `ifdef rtldump
      let clogpkt = rx_commitlog.u.first;
      rx_commitlog.u.deq;
      clogpkt.mode = csr.mv_prv;
			`ifdef hypervisor
				clogpkt.v = csr.mv_virtual;
			`endif
      rg_commitlog <= tagged Valid clogpkt;
    `endif
    end
    else begin
      `logLevel( stage5, 0, $format("[%2d]STAGE5 : Dropping instruction",hartid))
      wr_commit <= CommitData{addr: fuid.rd, data: ?, unlock_only:True
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu rdtype: fuid.rdtype `endif };
      rx_baseout.u.deq;
      rx_fuid.u.deq;
    `ifdef rtldump
      rx_commitlog.u.deq;
    `endif
    end
  endrule:rl_writeback_baseout

  /*doc:rule: This rule performs memory operations. In specific it completes a previously cached
  * store/atomic operation or initiates a new IO memory operation. This rule simply indicates the
  * Store buffer or the IO buffer held in the cache to initiate the respective operation. This
  * indication is basically a write to the wr_commit_cacheop/wr_commit_ioop wire with the current
  * epoch value.
  * In case a cached store/atomic op has to be dropped since the epochs don't match. The epoch value
  * sent will cause the respective entry in the caches to be dropped without any updates to cache/
  * memory*/
  rule rl_writeback_memop(rx_fuid.u.first.insttype == MEMORY );
    let memop = rx_memio.u.first;
    let fuid = rx_fuid.u.first;
    `logLevel( stage5, 0, $format("[%2d]STAGE5 : PC:%h",hartid,fuid.pc))
  `ifdef rtldump
    let clogpkt = rx_commitlog.u.first;
    CommitLogMem _pkt = ?;
    if (clogpkt.inst_type matches tagged MEM. cmem) 
      _pkt = cmem;
  `endif

    if (epochs_match) begin
    `ifdef dcache
      if (!memop.io) begin // cacheable store/atomic op
        `logLevel( stage5, 0, $format("[%2d]STAGE5 : Cached Store Op ",hartid, fshow(memop)))
        wr_commit_cacheop <= tuple2(rg_epoch, memop.sb_id);
        wr_increment_minstret <= True;
        rx_fuid.u.deq;
        rx_memio.u.deq;
      `ifdef atomic
        let cache_resp = memop.atomic_rd_data;
        if (memop.memaccess == Atomic) 
          wr_commit <= CommitData{addr: fuid.rd, data: zeroExtend(cache_resp), unlock_only:False
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu rdtype: fuid.rdtype `endif };
      `else
        Bit#(`elen) cache_resp = 0;
      `endif
      `ifdef rtldump
        rx_commitlog.u.deq;
        _pkt.commit_data = cache_resp;
        clogpkt.inst_type = tagged MEM _pkt;
        clogpkt.mode = csr.mv_prv;
			`ifdef hypervisor
				clogpkt.v = csr.mv_virtual;
			`endif
        rg_commitlog <= tagged Valid clogpkt;
      `endif
      end
      else 
    `endif
      begin 
        `logLevel( stage5, 0, $format("[%2d]STAGE5 : Non-Cached Memory Op ",hartid, fshow(memop)))
        if (!rg_ioop_init) begin
          rg_ioop_init <= True;
          wr_commit_ioop <= rg_epoch;
        end
        else if (wr_ioop_response matches tagged Valid .ioresp) begin
          rg_ioop_init <= False;
          if (ioresp.trap) begin
            let tvec <- csr.mav_upd_on_trap(ioresp.cause, fuid.pc, ioresp.word, ?);
            wr_flush <= WBFlush{flush: True, newpc : tvec, fencei: False 
                `ifdef supervisor , sfence: False `endif 
                `ifdef hypervisor , hfence: False `endif };
            `logLevel( stage5, 0, $format("[%2d]STAGE5 : Redirect PC:%h",hartid, tvec))
            rg_epoch <= ~rg_epoch;
            rx_fuid.u.deq;
            rx_memio.u.deq;
            wr_commit <= CommitData{addr: fuid.rd, data: ?, unlock_only: True
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu rdtype: fuid.rdtype `endif };
          `ifdef rtldump
            rx_commitlog.u.deq;
          `endif
          end
          else begin
            wr_increment_minstret <= True;
            let commit_data = ioresp.word;
            `ifdef spfpu if (memop.nanboxing) commit_data[63:32] = '1; `endif
            wr_commit <= CommitData{addr: fuid.rd, data: zeroExtend(commit_data), unlock_only:False
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu rdtype: fuid.rdtype `endif };
            rx_fuid.u.deq;
            rx_memio.u.deq;
          `ifdef rtldump
            rx_commitlog.u.deq;
            _pkt.commit_data = (fuid.rd ==0 `ifdef spfpu && fuid.rdtype == IRF `endif )?0:commit_data;
            clogpkt.inst_type = tagged MEM _pkt;
            clogpkt.mode = csr.mv_prv;
					`ifdef hypervisor
						clogpkt.v = csr.mv_virtual;
					`endif
            rg_commitlog <= tagged Valid clogpkt;
          `endif
          end
        end
        else begin
          `logLevel( stage5, 0, $format("[%2d]STAGE5: Waiting for IO response",hartid))
        end
      end
    end
    else begin
      `logLevel( stage5, 0, $format("[%2d]STAGE5 : Dropping instruction",hartid))
      wr_commit <= CommitData{addr: fuid.rd, data: ?, unlock_only:True
                                      `ifdef no_wawstalls , id: fuid.id `endif
                                      `ifdef spfpu rdtype: fuid.rdtype `endif };
      rx_memio.u.deq;
      rx_fuid.u.deq;
    `ifdef rtldump
      rx_commitlog.u.deq;
    `endif
    `ifdef dcache
      if(!memop.io)
        wr_commit_cacheop <= tuple2(rg_epoch, ?);
      else
    `endif
        wr_commit_ioop <= rg_epoch;
    end
  endrule:rl_writeback_memop

  /*doc:rule: This rule is fired when wr_increment_minstret is set and thus cases the minstret
  * register to increment*/
  rule rl_incr_minstret(wr_increment_minstret);
    csr.ma_incr_minstret(1);
  endrule:rl_incr_minstret

  interface rx = interface Ifc_s5_rx
    interface rx_systemout_from_stage4  = rx_systemout.e;
    interface rx_trapout_from_stage4  = rx_trapout.e;
    interface rx_baseout_from_stage4 = rx_baseout.e;
    interface rx_memio_from_stage4 = rx_memio.e;
    interface rx_fuid_from_stage4 = rx_fuid.e;
  `ifdef rtldump
    interface rx_commitlog = rx_commitlog.e;
  `endif
  endinterface;
  
  interface interrupts = interface Ifc_s5_interrupts
    method ma_clint_msip = csr.ma_set_mip_msip;
    method ma_clint_mtip = csr.ma_set_mip_mtip;
    method ma_clint_mtime = csr.ma_set_time;
    method ma_plic_meip = csr.ma_set_mip_meip;
  `ifdef hypervisor
  	method ma_plic_vseip = csr.ma_set_vseip;
  `endif
  `ifdef supervisor 
    method ma_plic_seip = csr.ma_set_mip_seip;
  `endif
  `ifdef usertraps
    method ma_plic_ueip = csr.ma_set_mip_ueip;
  `endif
  endinterface;
`ifdef debug 
  interface debug = interface Ifc_s5_debug
    method mv_csr_dcsr = csr.sbread.mv_csr_dcsr;
    method ma_debug_interrupt= csr.ma_set_mip_debug_interrupt;
    method mv_debug_mode= csr.mv_debug_mode;
    method mv_core_debugenable = csr.sbread.mv_csr_customcontrol[4];
    method mv_stop_timer = csr.mv_stop_timer;
    method mv_stop_count = csr.mv_stop_count;
  endinterface;
`endif

`ifdef perfmonitors
  interface perf = interface Ifc_s5_perfmonitors
    method ma_events = csr.ma_events;
   	method mv_count_exceptions = wr_count_exceptions;
   	method mv_count_interrupts = wr_count_interrupts;
   	method mv_count_csrops = wr_count_csrops;
   	method mv_count_microtraps = wr_count_microtrap;
  endinterface;
`endif
  
  interface common = interface Ifc_s5_common
    method mv_commit_rd = wr_commit;
    method mv_flush = wr_flush;
  `ifdef rtldump
    method mv_commit_log = rg_commitlog;
  `endif
  endinterface;
  
  interface cache = interface Ifc_s5_cache
    method mv_initiate_store = wr_commit_cacheop;
    method Bit#(1) mv_initiate_ioop = wr_commit_ioop;
    method Action ma_io_response(Maybe#(DMem_core_response#(TMul#(`dwords,8),`desize)) r);
      wr_ioop_response <= r;
    endmethod:ma_io_response
  endinterface;

  interface csrs = interface Ifc_s5_csrs;
    method mv_csr_misa_c = csr.sbread.mv_csr_misa[2];
    method mv_cacheenable = truncate(csr.sbread.mv_csr_customcontrol);
    method mv_curr_priv = pack(csr.mv_prv);
    method mv_csr_mstatus = csr.sbread.mv_csr_mstatus;
  `ifdef hypervisor
		`ifdef RV32
			method mv_csr_mstatush = csr.sbread.mv_csr_mstatush;
 		`endif
		method mv_csr_hstatus = csr.sbread.mv_csr_hstatus;
		method mv_csr_vsstatus = csr.sbread.mv_csr_vsstatus;				
		method mv_csr_vsatp = csr.sbread.mv_csr_vsatp;
		method mv_csr_hgatp = csr.sbread.mv_csr_hgatp;
		method mv_vs_bit = csr.mv_virtual;
  `endif
    method mv_csrs_to_decode = CSRtoDecode {prv: csr.mv_prv,
        csr_mip: truncate(csr.sbread.mv_csr_mip), 
        csr_mie: truncate(csr.sbread.mv_csr_mie), 
        csr_mstatus: truncate(csr.sbread.mv_csr_mstatus),
        csr_sstatus: `ifdef hypervisor (csr.mv_virtual == 1)? csr.sbread.mv_csr_vsstatus: `endif csr.sbread.mv_csr_mstatus,
        csr_misa: truncate(csr.sbread.mv_csr_misa)
      `ifdef spfpu
        ,frm: truncate(csr.sbread.mv_csr_frm)
      `endif
      `ifdef debug
        ,csr_dcsr: truncate(csr.sbread.mv_csr_dcsr)
      `endif
      `ifdef non_m_traps 
        ,csr_mideleg: truncate(csr.sbread.mv_csr_mideleg)
    `endif 
    `ifdef hypervisor
    , csr_hideleg: truncate(csr.sbread.mv_csr_hideleg)
    , csr_hstatus: truncate(csr.sbread.mv_csr_hstatus)   
    , csr_vs_bit: truncate(csr.mv_virtual)
      `endif };
    method mv_resume_wfi = unpack( |((csr.sbread.mv_csr_mip)& (csr.sbread.mv_csr_mie) ));
	`ifdef supervisor
		method mv_csr_satp = csr.sbread.mv_csr_satp;
	`endif
  `ifdef pmp
    method mv_pmp_cfg = csr.mv_pmpcfg;
    method mv_pmp_addr = csr.mv_pmpaddr;
  `endif
  `ifdef rtldump
    interface sbread = csr.sbread;
  `endif
  endinterface;
endmodule: mkstage5

endpackage: stage5

